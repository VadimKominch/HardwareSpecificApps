library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity counter_with_ts_signal is
  generic
  (
  Size:integer
  );
  port(
  reset:in std_logic;
  clk:in std_logic;
  Ts:out std_logic
  );
end counter_with_ts_signal;

architecture beh of counter_with_ts_signal is
signal count:std_logic_vector(Size-1 downto 0);
signal limit:std_logic_vector(Size-1 downto 0);

begin
  limit<=(others =>'1');
  process(clk)
    begin
      if(reset ='1') then
        count<=(others =>'0');
      elsif(rising_edge(clk)) then
        count<=count+1;
      end if;
    end process;
    --Comparison with max value
    Ts<='1' when count=limit else '0';
end beh;
