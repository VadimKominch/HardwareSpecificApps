library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;

entity addsub is
  generic(
  Size:integer);
  port(
  a:in std_logic_vector(Size-1 downto 0);
  b:in std_logic_vector(Size-1 downto 0);
  control:in std_logic;
  c:out std_logic_vector(Size-1 downto 0));
end addsub;

architecture beh of addsub is
begin
  process (a, b, control)
   begin 
   if control = '0' then 
   c <= a + b; 
   else 
   c <= a - b; 
   end if; 
  end process;
end beh;